module c432 (M1__PA, M2__PB, M3__PC, M5__Chan_3, M5__Chan_2, M5__Chan_1, 
    M5__Chan_0, E_8, E_7, E_6, E_5, E_4, E_3, E_2, E_1, E_0, A_8, A_7, A_6, A_5, 
    A_4, A_3, A_2, A_1, A_0, B_8, B_7, B_6, B_5, B_4, B_3, B_2, B_1, B_0, C_8, 
    C_7, C_6, C_5, C_4, C_3, C_2, C_1, C_0);

    input  E_8;
    input  E_7;
    input  E_6;
    input  E_5;
    input  E_4;
    input  E_3;
    input  E_2;
    input  E_1;
    input  E_0;
    input  A_8;
    input  A_7;
    input  A_6;
    input  A_5;
    input  A_4;
    input  A_3;
    input  A_2;
    input  A_1;
    input  A_0;
    input  B_8;
    input  B_7;
    input  B_6;
    input  B_5;
    input  B_4;
    input  B_3;
    input  B_2;
    input  B_1;
    input  B_0;
    input  C_8;
    input  C_7;
    input  C_6;
    input  C_5;
    input  C_4;
    input  C_3;
    input  C_2;
    input  C_1;
    input  C_0;

    output  M1__PA;
    output  M2__PB;
    output  M3__PC;
    output  M5__Chan_3;
    output  M5__Chan_2;
    output  M5__Chan_1;
    output  M5__Chan_0;

    inv1 M1__Ab0(.Y(M1__Ab_0), .A(A_0));
    inv1 M1__Ab1(.Y(M1__Ab_1), .A(A_1));
    inv1 M1__Ab2(.Y(M1__Ab_2), .A(A_2));
    inv1 M1__Ab3(.Y(M1__Ab_3), .A(A_3));
    inv1 M1__Ab4(.Y(M1__Ab_4), .A(A_4));
    inv1 M1__Ab5(.Y(M1__Ab_5), .A(A_5));
    inv1 M1__Ab6(.Y(M1__Ab_6), .A(A_6));
    inv1 M1__Ab7(.Y(M1__Ab_7), .A(A_7));
    inv1 M1__Ab8(.Y(M1__Ab_8), .A(A_8));
    nand2 M1__EAb0(.Y(M1__EAb_0), .A(M1__Ab_0), .B(E_0));
    nand2 M1__EAb1(.Y(M1__EAb_1), .A(M1__Ab_1), .B(E_1));
    nand2 M1__EAb2(.Y(M1__EAb_2), .A(M1__Ab_2), .B(E_2));
    nand2 M1__EAb3(.Y(M1__EAb_3), .A(M1__Ab_3), .B(E_3));
    nand2 M1__EAb4(.Y(M1__EAb_4), .A(M1__Ab_4), .B(E_4));
    nand2 M1__EAb5(.Y(M1__EAb_5), .A(M1__Ab_5), .B(E_5));
    nand2 M1__EAb6(.Y(M1__EAb_6), .A(M1__Ab_6), .B(E_6));
    nand2 M1__EAb7(.Y(M1__EAb_7), .A(M1__Ab_7), .B(E_7));
    nand2 M1__EAb8(.Y(M1__EAb_8), .A(M1__Ab_8), .B(E_8));
    nand2 M1__PAgate(.Y(M1__PA), .A(M1__PAi), .B(M1__EAb_8));
    and2 M1__PAigate(.Y(M1__PAi), .A(M1__PAi_2), .B(M1__PAi_t0));
    and2 M1__PAigate_0(.Y(M1__PAi_0), .A(M1__EAb_2), .B(M1__PAi_0_t0));
    and2 M1__PAigate_0_t0(.Y(M1__PAi_0_t0), .A(M1__EAb_0), .B(M1__EAb_1));
    and2 M1__PAigate_1(.Y(M1__PAi_1), .A(M1__EAb_5), .B(M1__PAi_1_t0));
    and2 M1__PAigate_1_t0(.Y(M1__PAi_1_t0), .A(M1__EAb_3), .B(M1__EAb_4));
    and2 M1__PAigate_2(.Y(M1__PAi_2), .A(M1__EAb_6), .B(M1__EAb_7));
    and2 M1__PAigate_t0(.Y(M1__PAi_t0), .A(M1__PAi_0), .B(M1__PAi_1));
    xor2 M1__X10(.Y(M1__X1_0), .A(M1__PA), .B(M1__EAb_0));
    xor2 M1__X11(.Y(M1__X1_1), .A(M1__PA), .B(M1__EAb_1));
    xor2 M1__X12(.Y(M1__X1_2), .A(M1__PA), .B(M1__EAb_2));
    xor2 M1__X13(.Y(M1__X1_3), .A(M1__PA), .B(M1__EAb_3));
    xor2 M1__X14(.Y(M1__X1_4), .A(M1__PA), .B(M1__EAb_4));
    xor2 M1__X15(.Y(M1__X1_5), .A(M1__PA), .B(M1__EAb_5));
    xor2 M1__X16(.Y(M1__X1_6), .A(M1__PA), .B(M1__EAb_6));
    xor2 M1__X17(.Y(M1__X1_7), .A(M1__PA), .B(M1__EAb_7));
    xor2 M1__X18(.Y(M1__X1_8), .A(M1__PA), .B(M1__EAb_8));
    inv1 M2__Eb0(.Y(M2__Eb_0), .A(E_0));
    inv1 M2__Eb1(.Y(M2__Eb_1), .A(E_1));
    inv1 M2__Eb2(.Y(M2__Eb_2), .A(E_2));
    inv1 M2__Eb3(.Y(M2__Eb_3), .A(E_3));
    inv1 M2__Eb4(.Y(M2__Eb_4), .A(E_4));
    inv1 M2__Eb5(.Y(M2__Eb_5), .A(E_5));
    inv1 M2__Eb6(.Y(M2__Eb_6), .A(E_6));
    inv1 M2__Eb7(.Y(M2__Eb_7), .A(E_7));
    inv1 M2__Eb8(.Y(M2__Eb_8), .A(E_8));
    nor2 M2__EbB0(.Y(M2__EbB_0), .A(M2__Eb_0), .B(B_0));
    nor2 M2__EbB1(.Y(M2__EbB_1), .A(M2__Eb_1), .B(B_1));
    nor2 M2__EbB2(.Y(M2__EbB_2), .A(M2__Eb_2), .B(B_2));
    nor2 M2__EbB3(.Y(M2__EbB_3), .A(M2__Eb_3), .B(B_3));
    nor2 M2__EbB4(.Y(M2__EbB_4), .A(M2__Eb_4), .B(B_4));
    nor2 M2__EbB5(.Y(M2__EbB_5), .A(M2__Eb_5), .B(B_5));
    nor2 M2__EbB6(.Y(M2__EbB_6), .A(M2__Eb_6), .B(B_6));
    nor2 M2__EbB7(.Y(M2__EbB_7), .A(M2__Eb_7), .B(B_7));
    nor2 M2__EbB8(.Y(M2__EbB_8), .A(M2__Eb_8), .B(B_8));
    nand2 M2__PBgate(.Y(M2__PB), .A(M2__PBi), .B(M2__XEB_8));
    and2 M2__PBigate(.Y(M2__PBi), .A(M2__PBi_2), .B(M2__PBi_t0));
    and2 M2__PBigate_0(.Y(M2__PBi_0), .A(M2__XEB_2), .B(M2__PBi_0_t0));
    and2 M2__PBigate_0_t0(.Y(M2__PBi_0_t0), .A(M2__XEB_0), .B(M2__XEB_1));
    and2 M2__PBigate_1(.Y(M2__PBi_1), .A(M2__XEB_5), .B(M2__PBi_1_t0));
    and2 M2__PBigate_1_t0(.Y(M2__PBi_1_t0), .A(M2__XEB_3), .B(M2__XEB_4));
    and2 M2__PBigate_2(.Y(M2__PBi_2), .A(M2__XEB_6), .B(M2__XEB_7));
    and2 M2__PBigate_t0(.Y(M2__PBi_t0), .A(M2__PBi_0), .B(M2__PBi_1));
    xor2 M2__X20(.Y(M2__X2_0), .A(M2__PB), .B(M2__XEB_0));
    xor2 M2__X21(.Y(M2__X2_1), .A(M2__PB), .B(M2__XEB_1));
    xor2 M2__X22(.Y(M2__X2_2), .A(M2__PB), .B(M2__XEB_2));
    xor2 M2__X23(.Y(M2__X2_3), .A(M2__PB), .B(M2__XEB_3));
    xor2 M2__X24(.Y(M2__X2_4), .A(M2__PB), .B(M2__XEB_4));
    xor2 M2__X25(.Y(M2__X2_5), .A(M2__PB), .B(M2__XEB_5));
    xor2 M2__X26(.Y(M2__X2_6), .A(M2__PB), .B(M2__XEB_6));
    xor2 M2__X27(.Y(M2__X2_7), .A(M2__PB), .B(M2__XEB_7));
    xor2 M2__X28(.Y(M2__X2_8), .A(M2__PB), .B(M2__XEB_8));
    nand2 M2__XEB0(.Y(M2__XEB_0), .A(M2__EbB_0), .B(M1__X1_0));
    nand2 M2__XEB1(.Y(M2__XEB_1), .A(M2__EbB_1), .B(M1__X1_1));
    nand2 M2__XEB2(.Y(M2__XEB_2), .A(M2__EbB_2), .B(M1__X1_2));
    nand2 M2__XEB3(.Y(M2__XEB_3), .A(M2__EbB_3), .B(M1__X1_3));
    nand2 M2__XEB4(.Y(M2__XEB_4), .A(M2__EbB_4), .B(M1__X1_4));
    nand2 M2__XEB5(.Y(M2__XEB_5), .A(M2__EbB_5), .B(M1__X1_5));
    nand2 M2__XEB6(.Y(M2__XEB_6), .A(M2__EbB_6), .B(M1__X1_6));
    nand2 M2__XEB7(.Y(M2__XEB_7), .A(M2__EbB_7), .B(M1__X1_7));
    nand2 M2__XEB8(.Y(M2__XEB_8), .A(M2__EbB_8), .B(M1__X1_8));
    inv1 M3__Eb0(.Y(M3__Eb_0), .A(E_0));
    inv1 M3__Eb1(.Y(M3__Eb_1), .A(E_1));
    inv1 M3__Eb2(.Y(M3__Eb_2), .A(E_2));
    inv1 M3__Eb3(.Y(M3__Eb_3), .A(E_3));
    inv1 M3__Eb4(.Y(M3__Eb_4), .A(E_4));
    inv1 M3__Eb5(.Y(M3__Eb_5), .A(E_5));
    inv1 M3__Eb6(.Y(M3__Eb_6), .A(E_6));
    inv1 M3__Eb7(.Y(M3__Eb_7), .A(E_7));
    inv1 M3__Eb8(.Y(M3__Eb_8), .A(E_8));
    nor2 M3__EbC0(.Y(M3__EbC_0), .A(M3__Eb_0), .B(C_0));
    nor2 M3__EbC1(.Y(M3__EbC_1), .A(M3__Eb_1), .B(C_1));
    nor2 M3__EbC2(.Y(M3__EbC_2), .A(M3__Eb_2), .B(C_2));
    nor2 M3__EbC3(.Y(M3__EbC_3), .A(M3__Eb_3), .B(C_3));
    nor2 M3__EbC4(.Y(M3__EbC_4), .A(M3__Eb_4), .B(C_4));
    nor2 M3__EbC5(.Y(M3__EbC_5), .A(M3__Eb_5), .B(C_5));
    nor2 M3__EbC6(.Y(M3__EbC_6), .A(M3__Eb_6), .B(C_6));
    nor2 M3__EbC7(.Y(M3__EbC_7), .A(M3__Eb_7), .B(C_7));
    nor2 M3__EbC8(.Y(M3__EbC_8), .A(M3__Eb_8), .B(C_8));
    nand2 M3__PCgate(.Y(M3__PC), .A(M3__PCi), .B(M3__XEC_8));
    and2 M3__PCigate(.Y(M3__PCi), .A(M3__PCi_2), .B(M3__PCi_t0));
    and2 M3__PCigate_0(.Y(M3__PCi_0), .A(M3__XEC_2), .B(M3__PCi_0_t0));
    and2 M3__PCigate_0_t0(.Y(M3__PCi_0_t0), .A(M3__XEC_0), .B(M3__XEC_1));
    and2 M3__PCigate_1(.Y(M3__PCi_1), .A(M3__XEC_5), .B(M3__PCi_1_t0));
    and2 M3__PCigate_1_t0(.Y(M3__PCi_1_t0), .A(M3__XEC_3), .B(M3__XEC_4));
    and2 M3__PCigate_2(.Y(M3__PCi_2), .A(M3__XEC_6), .B(M3__XEC_7));
    and2 M3__PCigate_t0(.Y(M3__PCi_t0), .A(M3__PCi_0), .B(M3__PCi_1));
    nand2 M3__XEC0(.Y(M3__XEC_0), .A(M2__X2_0), .B(M3__XEC_0_t0));
    and2 M3__XEC0_t0(.Y(M3__XEC_0_t0), .A(M3__EbC_0), .B(M1__X1_0));
    nand2 M3__XEC1(.Y(M3__XEC_1), .A(M2__X2_1), .B(M3__XEC_1_t0));
    and2 M3__XEC1_t0(.Y(M3__XEC_1_t0), .A(M3__EbC_1), .B(M1__X1_1));
    nand2 M3__XEC2(.Y(M3__XEC_2), .A(M2__X2_2), .B(M3__XEC_2_t0));
    and2 M3__XEC2_t0(.Y(M3__XEC_2_t0), .A(M3__EbC_2), .B(M1__X1_2));
    nand2 M3__XEC3(.Y(M3__XEC_3), .A(M2__X2_3), .B(M3__XEC_3_t0));
    and2 M3__XEC3_t0(.Y(M3__XEC_3_t0), .A(M3__EbC_3), .B(M1__X1_3));
    nand2 M3__XEC4(.Y(M3__XEC_4), .A(M2__X2_4), .B(M3__XEC_4_t0));
    and2 M3__XEC4_t0(.Y(M3__XEC_4_t0), .A(M3__EbC_4), .B(M1__X1_4));
    nand2 M3__XEC5(.Y(M3__XEC_5), .A(M2__X2_5), .B(M3__XEC_5_t0));
    and2 M3__XEC5_t0(.Y(M3__XEC_5_t0), .A(M3__EbC_5), .B(M1__X1_5));
    nand2 M3__XEC6(.Y(M3__XEC_6), .A(M2__X2_6), .B(M3__XEC_6_t0));
    and2 M3__XEC6_t0(.Y(M3__XEC_6_t0), .A(M3__EbC_6), .B(M1__X1_6));
    nand2 M3__XEC7(.Y(M3__XEC_7), .A(M2__X2_7), .B(M3__XEC_7_t0));
    and2 M3__XEC7_t0(.Y(M3__XEC_7_t0), .A(M3__EbC_7), .B(M1__X1_7));
    nand2 M3__XEC8(.Y(M3__XEC_8), .A(M2__X2_8), .B(M3__XEC_8_t0));
    and2 M3__XEC8_t0(.Y(M3__XEC_8_t0), .A(M3__EbC_8), .B(M1__X1_8));
    nand2 M4__APA0(.Y(M4__APA_0), .A(A_0), .B(M1__PA));
    nand2 M4__APA1(.Y(M4__APA_1), .A(A_1), .B(M1__PA));
    nand2 M4__APA2(.Y(M4__APA_2), .A(A_2), .B(M1__PA));
    nand2 M4__APA3(.Y(M4__APA_3), .A(A_3), .B(M1__PA));
    nand2 M4__APA4(.Y(M4__APA_4), .A(A_4), .B(M1__PA));
    nand2 M4__APA5(.Y(M4__APA_5), .A(A_5), .B(M1__PA));
    nand2 M4__APA6(.Y(M4__APA_6), .A(A_6), .B(M1__PA));
    nand2 M4__APA7(.Y(M4__APA_7), .A(A_7), .B(M1__PA));
    nand2 M4__APA8(.Y(M4__APA_8), .A(A_8), .B(M1__PA));
    nand2 M4__BPB0(.Y(M4__BPB_0), .A(B_0), .B(M2__PB));
    nand2 M4__BPB1(.Y(M4__BPB_1), .A(B_1), .B(M2__PB));
    nand2 M4__BPB2(.Y(M4__BPB_2), .A(B_2), .B(M2__PB));
    nand2 M4__BPB3(.Y(M4__BPB_3), .A(B_3), .B(M2__PB));
    nand2 M4__BPB4(.Y(M4__BPB_4), .A(B_4), .B(M2__PB));
    nand2 M4__BPB5(.Y(M4__BPB_5), .A(B_5), .B(M2__PB));
    nand2 M4__BPB6(.Y(M4__BPB_6), .A(B_6), .B(M2__PB));
    nand2 M4__BPB7(.Y(M4__BPB_7), .A(B_7), .B(M2__PB));
    nand2 M4__BPB8(.Y(M4__BPB_8), .A(B_8), .B(M2__PB));
    nand2 M4__CPC0(.Y(M4__CPC_0), .A(C_0), .B(M3__PC));
    nand2 M4__CPC1(.Y(M4__CPC_1), .A(C_1), .B(M3__PC));
    nand2 M4__CPC2(.Y(M4__CPC_2), .A(C_2), .B(M3__PC));
    nand2 M4__CPC3(.Y(M4__CPC_3), .A(C_3), .B(M3__PC));
    nand2 M4__CPC4(.Y(M4__CPC_4), .A(C_4), .B(M3__PC));
    nand2 M4__CPC5(.Y(M4__CPC_5), .A(C_5), .B(M3__PC));
    nand2 M4__CPC6(.Y(M4__CPC_6), .A(C_6), .B(M3__PC));
    nand2 M4__CPC7(.Y(M4__CPC_7), .A(C_7), .B(M3__PC));
    nand2 M4__CPC8(.Y(M4__CPC_8), .A(C_8), .B(M3__PC));
    nand2 M4__I0(.Y(M4__I_0), .A(M4__I_0_t0), .B(M4__I_0_t1));
    and2 M4__I0_t0(.Y(M4__I_0_t0), .A(E_0), .B(M4__APA_0));
    and2 M4__I0_t1(.Y(M4__I_0_t1), .A(M4__BPB_0), .B(M4__CPC_0));
    nand2 M4__I1(.Y(M4__I_1), .A(M4__I_1_t0), .B(M4__I_1_t1));
    and2 M4__I1_t0(.Y(M4__I_1_t0), .A(E_1), .B(M4__APA_1));
    and2 M4__I1_t1(.Y(M4__I_1_t1), .A(M4__BPB_1), .B(M4__CPC_1));
    nand2 M4__I2(.Y(M4__I_2), .A(M4__I_2_t0), .B(M4__I_2_t1));
    and2 M4__I2_t0(.Y(M4__I_2_t0), .A(E_2), .B(M4__APA_2));
    and2 M4__I2_t1(.Y(M4__I_2_t1), .A(M4__BPB_2), .B(M4__CPC_2));
    nand2 M4__I3(.Y(M4__I_3), .A(M4__I_3_t0), .B(M4__I_3_t1));
    and2 M4__I3_t0(.Y(M4__I_3_t0), .A(E_3), .B(M4__APA_3));
    and2 M4__I3_t1(.Y(M4__I_3_t1), .A(M4__BPB_3), .B(M4__CPC_3));
    nand2 M4__I4(.Y(M4__I_4), .A(M4__I_4_t0), .B(M4__I_4_t1));
    and2 M4__I4_t0(.Y(M4__I_4_t0), .A(E_4), .B(M4__APA_4));
    and2 M4__I4_t1(.Y(M4__I_4_t1), .A(M4__BPB_4), .B(M4__CPC_4));
    nand2 M4__I5(.Y(M4__I_5), .A(M4__I_5_t0), .B(M4__I_5_t1));
    and2 M4__I5_t0(.Y(M4__I_5_t0), .A(E_5), .B(M4__APA_5));
    and2 M4__I5_t1(.Y(M4__I_5_t1), .A(M4__BPB_5), .B(M4__CPC_5));
    nand2 M4__I6(.Y(M4__I_6), .A(M4__I_6_t0), .B(M4__I_6_t1));
    and2 M4__I6_t0(.Y(M4__I_6_t0), .A(E_6), .B(M4__APA_6));
    and2 M4__I6_t1(.Y(M4__I_6_t1), .A(M4__BPB_6), .B(M4__CPC_6));
    nand2 M4__I7(.Y(M4__I_7), .A(M4__I_7_t0), .B(M4__I_7_t1));
    and2 M4__I7_t0(.Y(M4__I_7_t0), .A(E_7), .B(M4__APA_7));
    and2 M4__I7_t1(.Y(M4__I_7_t1), .A(M4__BPB_7), .B(M4__CPC_7));
    nand2 M4__I8(.Y(M4__I_8), .A(M4__I_8_t0), .B(M4__I_8_t1));
    and2 M4__I8_t0(.Y(M4__I_8_t0), .A(E_8), .B(M4__APA_8));
    and2 M4__I8_t1(.Y(M4__I_8_t1), .A(M4__BPB_8), .B(M4__CPC_8));
    nand2 M5__Chan0(.Y(M5__Chan_0), .A(M5__Chan_0_t0), .B(M5__Chan_0_t1));
    and2 M5__Chan0_t0(.Y(M5__Chan_0_t0), .A(M4__I_7), .B(M5__I56));
    and2 M5__Chan0_t1(.Y(M5__Chan_0_t1), .A(M5__I1256), .B(M5__I3456));
    nand2 M5__Chan1(.Y(M5__Chan_1), .A(M5__Chan_1_t0), .B(M5__Chan_1_t1));
    and2 M5__Chan1_t0(.Y(M5__Chan_1_t0), .A(M4__I_6), .B(M4__I_7));
    and2 M5__Chan1_t1(.Y(M5__Chan_1_t1), .A(M5__I245), .B(M5__I3456));
    nand2 M5__Chan2(.Y(M5__Chan_2), .A(M5__Chan_2_t0), .B(M5__Chan_2_t1));
    and2 M5__Chan2_t0(.Y(M5__Chan_2_t0), .A(M4__I_4), .B(M4__I_6));
    and2 M5__Chan2_t1(.Y(M5__Chan_2_t1), .A(M4__I_7), .B(M5__I56));
    nor2 M5__Chan3(.Y(M5__Chan_3), .A(M5__Iand), .B(M5__Ib8));
    nand2 M5__I1256gate(.Y(M5__I1256), .A(M5__I1256_t0), .B(M5__I1256_t1));
    and2 M5__I1256gate_t0(.Y(M5__I1256_t0), .A(M5__Ib1), .B(M4__I_2));
    and2 M5__I1256gate_t1(.Y(M5__I1256_t1), .A(M4__I_5), .B(M4__I_6));
    nand2 M5__I245gate(.Y(M5__I245), .A(M4__I_5), .B(M5__I245_t0));
    and2 M5__I245gate_t0(.Y(M5__I245_t0), .A(M5__Ib2), .B(M4__I_4));
    nand2 M5__I3456gate(.Y(M5__I3456), .A(M5__I3456_t0), .B(M5__I3456_t1));
    and2 M5__I3456gate_t0(.Y(M5__I3456_t0), .A(M5__Ib3), .B(M4__I_4));
    and2 M5__I3456gate_t1(.Y(M5__I3456_t1), .A(M4__I_5), .B(M4__I_6));
    nand2 M5__I56gate(.Y(M5__I56), .A(M5__Ib5), .B(M4__I_6));
    and2 M5__Iandgate(.Y(M5__Iand), .A(M5__Iand_2), .B(M5__Iand_t0));
    and2 M5__Iandgate_0(.Y(M5__Iand_0), .A(M4__I_2), .B(M5__Iand_0_t0));
    and2 M5__Iandgate_0_t0(.Y(M5__Iand_0_t0), .A(M4__I_0), .B(M4__I_1));
    and2 M5__Iandgate_1(.Y(M5__Iand_1), .A(M4__I_5), .B(M5__Iand_1_t0));
    and2 M5__Iandgate_1_t0(.Y(M5__Iand_1_t0), .A(M4__I_3), .B(M4__I_4));
    and2 M5__Iandgate_2(.Y(M5__Iand_2), .A(M4__I_6), .B(M4__I_7));
    and2 M5__Iandgate_t0(.Y(M5__Iand_t0), .A(M5__Iand_0), .B(M5__Iand_1));
    inv1 M5__Ib1gate(.Y(M5__Ib1), .A(M4__I_1));
    inv1 M5__Ib2gate(.Y(M5__Ib2), .A(M4__I_2));
    inv1 M5__Ib3gate(.Y(M5__Ib3), .A(M4__I_3));
    inv1 M5__Ib5gate(.Y(M5__Ib5), .A(M4__I_5));
    inv1 M5__Ib8gate(.Y(M5__Ib8), .A(M4__I_8));

endmodule /* c432 */

